// erro
